`ifndef __TEST_TOP_SVH__
`define __TEST_TOP_SVH__

`include "base_test.svh"
`include "order_data_multi_test.svh"
`include "random_data_multi_test.svh"
`include "input_always_valid_test.svh"

`endif
